module sdram (
	clk,
	rst
);

input clk;
input rst;


endmodule 
