//top.v

/**
 * Used as a staging area for demoing all the design.
 *	Demonstrates the following code
 *		<??>_io_handler
 *		wishbone_master
 *		wishbone_interconnect
 *		wishbone_rom
 *		wishbone_slave
 *
 */

module top (
	clk,
	rst	
);

input clk;
input rst;

endmodule
