//dot_tb.v

module dot_tb (
);


endmodule
